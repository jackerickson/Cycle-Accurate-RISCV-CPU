module counter
    (
        input [3:0] x,
        output [3:0] z
    );
    assign z = x + 1;

endmodule // counter
